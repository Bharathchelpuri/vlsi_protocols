program apb_test;
apb_env env_h;

initial begin 
env_h=new();
env_h.env_main();
end 

endprogram 
